module hello (
    hello
);
    
endmodule