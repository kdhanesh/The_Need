module uart_rtl (
    
);
    
endmodule